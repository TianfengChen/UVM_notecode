typedef uvm_sequence #(transact) my_sequencer;